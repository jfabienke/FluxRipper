//==============================================================================
// ISA Plug-and-Play Controller
//==============================================================================
// File: isa_pnp_controller.v
// Description: ISA PnP protocol implementation for automatic resource
//              configuration. Supports both FDC and WD HDD controllers.
//
// Features:
//   - PnP initiation key detection (32-byte sequence)
//   - Serial isolation protocol
//   - Two logical devices: FDC (LD0) and WD (LD1)
//   - Dynamic I/O base and IRQ configuration
//   - Resource descriptor ROM
//   - Integration with isa_pnp_sniffer for "Sleep-until-Key" strategy
//   - Legacy mode support for non-PnP systems
//
// PnP Port Map:
//   0x279 - Address port (write-only)
//   0xA79 - Write Data port
//   0x20B - Read Data port (configurable)
//
// Integration with Auto-Config:
//   - Sniffer detects initiation key and signals pnp_key_valid
//   - Controller starts in ST_WAIT_KEY but legacy I/O remains active
//   - Upon key detection, transitions to ST_ISOLATION
//   - Returns to legacy mode via CC_WAIT_FOR_KEY command
//
// Author: Claude Code (FluxRipper Project)
// Date: 2025-12-04 21:55
// Updated: 2025-12-07 - Added sniffer integration for universal compatibility
//==============================================================================

`timescale 1ns / 1ps

module isa_pnp_controller #(
    // EISA Vendor ID: "FLX" encoded (0x0C1F = F, L, X compressed)
    parameter [31:0] VENDOR_ID = 32'h0C1F1234,
    // Device serial number
    parameter [31:0] SERIAL_NUM = 32'h00000001
)(
    input  wire        clk,
    input  wire        reset_n,

    //=========================================================================
    // ISA Bus Interface
    //=========================================================================
    input  wire [9:0]  isa_addr,
    input  wire [7:0]  isa_data_in,
    output reg  [7:0]  isa_data_out,
    output wire        isa_data_oe,
    input  wire        isa_ior_n,
    input  wire        isa_iow_n,
    input  wire        isa_aen,

    //=========================================================================
    // Configured Resources (outputs to address decoder)
    //=========================================================================
    // FDC Configuration (Logical Device 0)
    output reg         fdc_activated,
    output reg  [9:0]  fdc_io_base,        // Default 0x3F0
    output reg  [3:0]  fdc_irq,            // Default IRQ6
    output reg  [2:0]  fdc_dma,            // Default DRQ2

    // WD Configuration (Logical Device 1)
    output reg         wd_activated,
    output reg  [9:0]  wd_io_base,         // Default 0x1F0
    output reg  [9:0]  wd_alt_base,        // Default 0x3F6
    output reg  [3:0]  wd_irq,             // Default IRQ14 (AT) / IRQ5 (XT)
    output reg  [2:0]  wd_dma,             // Default DRQ3 (XT mode)

    //=========================================================================
    // Status
    //=========================================================================
    output reg         pnp_configured,     // PnP configuration complete
    output reg  [7:0]  pnp_csn,            // Assigned Card Select Number

    //=========================================================================
    // Auto-Config Integration (Sniffer Interface)
    //=========================================================================
    input  wire        pnp_key_valid,      // Sniffer detected valid initiation key
    input  wire        legacy_mode_req,    // Request return to legacy mode
    output wire        pnp_config_active,  // In PnP configuration mode
    output wire        return_to_legacy    // Signal return to Wait-for-Key
);

    //=========================================================================
    // PnP Protocol Constants
    //=========================================================================
    localparam ADDR_PORT     = 10'h279;
    localparam WRITE_PORT    = 10'hA79;
    localparam READ_PORT_DEF = 10'h20B;    // Default read data port

    // PnP Register Addresses
    localparam REG_SET_RD_DATA   = 8'h00;
    localparam REG_SERIAL_ISOL   = 8'h01;
    localparam REG_CONFIG_CTRL   = 8'h02;
    localparam REG_WAKE          = 8'h03;
    localparam REG_RESOURCE_DATA = 8'h04;
    localparam REG_STATUS        = 8'h05;
    localparam REG_CSN           = 8'h06;
    localparam REG_LOG_DEV       = 8'h07;

    // Logical Device Registers (base + offset)
    localparam REG_ACTIVATE      = 8'h30;
    localparam REG_IO_RANGE_CHK  = 8'h31;
    localparam REG_IO_BASE_HI    = 8'h60;
    localparam REG_IO_BASE_LO    = 8'h61;
    localparam REG_IO2_BASE_HI   = 8'h62;
    localparam REG_IO2_BASE_LO   = 8'h63;
    localparam REG_IRQ_SELECT    = 8'h70;
    localparam REG_IRQ_TYPE      = 8'h71;
    localparam REG_DMA_SELECT    = 8'h74;

    // Config Control bits
    localparam CC_RESET          = 8'h01;
    localparam CC_WAIT_FOR_KEY   = 8'h02;
    localparam CC_RETURN_CSN     = 8'h04;

    //=========================================================================
    // PnP Initiation Key (LFSR sequence)
    //=========================================================================
    // The 32-byte initiation key is generated by an LFSR
    // Starting value: 0x6A, polynomial: x^8 + x^4 + x^3 + x^2 + 1

    reg [7:0] key_lfsr;
    reg [4:0] key_count;
    wire key_match = (key_count == 5'd32);

    wire [7:0] lfsr_next = {key_lfsr[6:0],
                           key_lfsr[7] ^ key_lfsr[3] ^ key_lfsr[2] ^ key_lfsr[1]};

    //=========================================================================
    // State Machine
    //=========================================================================
    localparam [3:0] ST_WAIT_KEY   = 4'd0;   // Waiting for initiation key
    localparam [3:0] ST_ISOLATION  = 4'd1;   // Serial isolation protocol
    localparam [3:0] ST_CONFIG     = 4'd2;   // Configuration mode
    localparam [3:0] ST_SLEEP      = 4'd3;   // Sleep state

    reg [3:0] state;

    //=========================================================================
    // Internal Registers
    //=========================================================================
    reg [7:0]  current_addr;       // Current register address
    reg [7:0]  current_ld;         // Current logical device
    reg [9:0]  read_data_port;     // Configured read data port
    reg [7:0]  isolation_byte;     // Current byte in isolation
    reg [2:0]  isolation_bit;      // Current bit in isolation
    reg        isolation_active;   // In isolation sequence

    // Resource data ROM pointer
    reg [7:0]  resource_ptr;
    reg        resource_ready;

    // Return to legacy mode signal
    reg        return_legacy_r;

    //=========================================================================
    // ISA Port Decoding
    //=========================================================================
    wire addr_port_sel  = (isa_addr == ADDR_PORT) && !isa_aen;
    wire write_port_sel = (isa_addr == WRITE_PORT) && !isa_aen;
    wire read_port_sel  = (isa_addr == read_data_port) && !isa_aen;

    // Edge detection
    reg isa_iow_n_d;
    wire write_strobe = isa_iow_n_d && !isa_iow_n;

    always @(posedge clk) begin
        isa_iow_n_d <= isa_iow_n;
    end

    //=========================================================================
    // Resource Data ROM
    //=========================================================================
    // Contains PnP resource descriptors for FDC and WD

    wire [7:0] resource_data;

    isa_pnp_rom #(
        .VENDOR_ID(VENDOR_ID),
        .SERIAL_NUM(SERIAL_NUM)
    ) u_resource_rom (
        .clk(clk),
        .addr(resource_ptr),
        .data(resource_data)
    );

    //=========================================================================
    // Main State Machine
    //=========================================================================
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            state            <= ST_WAIT_KEY;
            current_addr     <= 8'h00;
            current_ld       <= 8'h00;
            read_data_port   <= READ_PORT_DEF;
            pnp_csn          <= 8'h00;
            pnp_configured   <= 1'b0;

            // Default FDC configuration
            fdc_activated    <= 1'b0;
            fdc_io_base      <= 10'h3F0;
            fdc_irq          <= 4'd6;
            fdc_dma          <= 3'd2;

            // Default WD configuration
            wd_activated     <= 1'b0;
            wd_io_base       <= 10'h1F0;
            wd_alt_base      <= 10'h3F6;
            wd_irq           <= 4'd14;
            wd_dma           <= 3'd3;     // DRQ3 for XT mode

            // Key detection
            key_lfsr         <= 8'h6A;
            key_count        <= 5'd0;

            // Isolation
            isolation_byte   <= 8'h00;
            isolation_bit    <= 3'd0;
            isolation_active <= 1'b0;

            // Resource ROM
            resource_ptr     <= 8'h00;
            resource_ready   <= 1'b0;

            // Legacy return signal
            return_legacy_r  <= 1'b0;

        end else begin
            // Handle sniffer key detection (external trigger)
            if (pnp_key_valid && state == ST_WAIT_KEY) begin
                // Sniffer has validated the 32-byte key
                // Transition directly to isolation mode
                state     <= ST_ISOLATION;
                key_count <= 5'd0;
                key_lfsr  <= 8'h6A;
            end

            // Handle external legacy mode request
            if (legacy_mode_req) begin
                state           <= ST_WAIT_KEY;
                return_legacy_r <= 1'b1;
            end else begin
                return_legacy_r <= 1'b0;
            end
            // Default: clear one-shot signals
            resource_ready <= 1'b0;

            case (state)
                //-------------------------------------------------------------
                ST_WAIT_KEY: begin
                    // Wait for 32-byte initiation key
                    // NOTE: With sniffer integration, key detection is handled by
                    // isa_pnp_sniffer.v which validates the key and sets pnp_key_valid.
                    // This internal key detection is kept as fallback/redundancy.
                    //
                    // IMPORTANT: While in ST_WAIT_KEY, the card remains ACTIVE in
                    // legacy mode - responding to default I/O addresses (0x3F0, 0x1F0).
                    // This ensures compatibility with non-PnP systems.

                    if (write_strobe && addr_port_sel) begin
                        if (isa_data_in == key_lfsr) begin
                            key_count <= key_count + 1'b1;
                            key_lfsr  <= lfsr_next;

                            if (key_count == 5'd31) begin
                                // Key complete - enter isolation
                                state     <= ST_ISOLATION;
                                key_count <= 5'd0;
                                key_lfsr  <= 8'h6A;
                            end
                        end else begin
                            // Mismatch - reset key detection
                            key_count <= 5'd0;
                            key_lfsr  <= 8'h6A;
                        end
                    end
                end

                //-------------------------------------------------------------
                ST_ISOLATION: begin
                    // Serial isolation protocol
                    if (write_strobe && addr_port_sel) begin
                        current_addr <= isa_data_in;

                        // Handle isolation commands
                        if (isa_data_in == REG_SERIAL_ISOL) begin
                            // Start isolation sequence
                            isolation_active <= 1'b1;
                            isolation_byte   <= VENDOR_ID[7:0];  // First byte
                            isolation_bit    <= 3'd0;
                        end else if (isa_data_in == REG_CONFIG_CTRL) begin
                            // Will handle in write port
                        end else if (isa_data_in == REG_CSN) begin
                            // CSN assignment
                        end else if (isa_data_in == REG_WAKE) begin
                            // Wake command
                        end
                    end

                    if (write_strobe && write_port_sel) begin
                        case (current_addr)
                            REG_SET_RD_DATA: begin
                                // Set read data port address
                                read_data_port <= {2'b00, isa_data_in};
                            end

                            REG_CONFIG_CTRL: begin
                                if (isa_data_in & CC_RESET) begin
                                    state <= ST_WAIT_KEY;
                                end
                                if (isa_data_in & CC_WAIT_FOR_KEY) begin
                                    state <= ST_WAIT_KEY;
                                end
                            end

                            REG_CSN: begin
                                // Assign Card Select Number
                                pnp_csn <= isa_data_in;
                                if (isa_data_in != 8'h00) begin
                                    state          <= ST_CONFIG;
                                    pnp_configured <= 1'b1;
                                end
                            end

                            REG_WAKE: begin
                                // Wake card with specific CSN
                                if (isa_data_in == pnp_csn && pnp_csn != 8'h00) begin
                                    state <= ST_CONFIG;
                                end
                            end
                        endcase
                    end
                end

                //-------------------------------------------------------------
                ST_CONFIG: begin
                    // Configuration mode - handle logical device configuration
                    if (write_strobe && addr_port_sel) begin
                        current_addr <= isa_data_in;
                    end

                    if (write_strobe && write_port_sel) begin
                        case (current_addr)
                            REG_CONFIG_CTRL: begin
                                if (isa_data_in & CC_WAIT_FOR_KEY) begin
                                    state <= ST_WAIT_KEY;
                                end
                            end

                            REG_WAKE: begin
                                // Re-enter config for specific CSN
                                if (isa_data_in == pnp_csn) begin
                                    // Already in config
                                end else if (isa_data_in == 8'h00) begin
                                    state <= ST_ISOLATION;
                                end
                            end

                            REG_LOG_DEV: begin
                                // Select logical device
                                current_ld <= isa_data_in;
                            end

                            REG_ACTIVATE: begin
                                // Activate/deactivate logical device
                                if (current_ld == 8'h00) begin
                                    fdc_activated <= (isa_data_in & 8'h01) != 0;
                                end else if (current_ld == 8'h01) begin
                                    wd_activated <= (isa_data_in & 8'h01) != 0;
                                end
                            end

                            REG_IO_BASE_HI: begin
                                if (current_ld == 8'h00) begin
                                    fdc_io_base[9:8] <= isa_data_in[1:0];
                                end else if (current_ld == 8'h01) begin
                                    wd_io_base[9:8] <= isa_data_in[1:0];
                                end
                            end

                            REG_IO_BASE_LO: begin
                                if (current_ld == 8'h00) begin
                                    fdc_io_base[7:0] <= isa_data_in;
                                end else if (current_ld == 8'h01) begin
                                    wd_io_base[7:0] <= isa_data_in;
                                end
                            end

                            REG_IO2_BASE_HI: begin
                                // Secondary I/O base (WD alternate)
                                if (current_ld == 8'h01) begin
                                    wd_alt_base[9:8] <= isa_data_in[1:0];
                                end
                            end

                            REG_IO2_BASE_LO: begin
                                if (current_ld == 8'h01) begin
                                    wd_alt_base[7:0] <= isa_data_in;
                                end
                            end

                            REG_IRQ_SELECT: begin
                                if (current_ld == 8'h00) begin
                                    fdc_irq <= isa_data_in[3:0];
                                end else if (current_ld == 8'h01) begin
                                    wd_irq <= isa_data_in[3:0];
                                end
                            end

                            REG_DMA_SELECT: begin
                                if (current_ld == 8'h00) begin
                                    fdc_dma <= isa_data_in[2:0];
                                end else if (current_ld == 8'h01) begin
                                    wd_dma <= isa_data_in[2:0];
                                end
                            end
                        endcase
                    end
                end

                //-------------------------------------------------------------
                ST_SLEEP: begin
                    // Sleep state - only respond to wake commands
                    if (write_strobe && addr_port_sel && isa_data_in == REG_WAKE) begin
                        // Will check CSN in write port
                    end

                    if (write_strobe && write_port_sel && current_addr == REG_WAKE) begin
                        if (isa_data_in == pnp_csn) begin
                            state <= ST_CONFIG;
                        end
                    end
                end

                //-------------------------------------------------------------
                default: begin
                    state <= ST_WAIT_KEY;
                end
            endcase
        end
    end

    //=========================================================================
    // Read Data Output
    //=========================================================================
    always @(*) begin
        isa_data_out = 8'hFF;

        if (read_port_sel && !isa_ior_n) begin
            case (current_addr)
                REG_SERIAL_ISOL: begin
                    // Return isolation bit (duplicated)
                    if (isolation_active) begin
                        isa_data_out = isolation_byte[isolation_bit] ?
                                       8'h55 : 8'hAA;
                    end
                end

                REG_RESOURCE_DATA: begin
                    // Return resource ROM data
                    isa_data_out = resource_data;
                end

                REG_STATUS: begin
                    // Resource data status
                    isa_data_out = resource_ready ? 8'h01 : 8'h00;
                end

                REG_CSN: begin
                    isa_data_out = pnp_csn;
                end

                REG_LOG_DEV: begin
                    isa_data_out = current_ld;
                end

                REG_ACTIVATE: begin
                    if (current_ld == 8'h00) begin
                        isa_data_out = {7'b0, fdc_activated};
                    end else if (current_ld == 8'h01) begin
                        isa_data_out = {7'b0, wd_activated};
                    end
                end

                REG_IO_BASE_HI: begin
                    if (current_ld == 8'h00) begin
                        isa_data_out = {6'b0, fdc_io_base[9:8]};
                    end else if (current_ld == 8'h01) begin
                        isa_data_out = {6'b0, wd_io_base[9:8]};
                    end
                end

                REG_IO_BASE_LO: begin
                    if (current_ld == 8'h00) begin
                        isa_data_out = fdc_io_base[7:0];
                    end else if (current_ld == 8'h01) begin
                        isa_data_out = wd_io_base[7:0];
                    end
                end

                REG_IRQ_SELECT: begin
                    if (current_ld == 8'h00) begin
                        isa_data_out = {4'b0, fdc_irq};
                    end else if (current_ld == 8'h01) begin
                        isa_data_out = {4'b0, wd_irq};
                    end
                end

                REG_DMA_SELECT: begin
                    if (current_ld == 8'h00) begin
                        isa_data_out = {5'b0, fdc_dma};
                    end else if (current_ld == 8'h01) begin
                        isa_data_out = {5'b0, wd_dma};
                    end else begin
                        isa_data_out = 8'h04;  // No DMA (value 4)
                    end
                end

                default: begin
                    isa_data_out = 8'hFF;
                end
            endcase
        end
    end

    // Output enable for read data port
    assign isa_data_oe = read_port_sel && !isa_ior_n && !isa_aen &&
                         (state == ST_ISOLATION || state == ST_CONFIG);

    //=========================================================================
    // Auto-Config Status Outputs
    //=========================================================================
    // PnP configuration mode active (isolation or config states)
    assign pnp_config_active = (state == ST_ISOLATION) || (state == ST_CONFIG);

    // Signal to sniffer/auto-config that we've returned to wait-for-key
    assign return_to_legacy = return_legacy_r || (state == ST_WAIT_KEY && !pnp_key_valid);

endmodule
